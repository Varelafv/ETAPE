----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 28.09.2022 16:47:14
-- Design Name: 
-- Module Name: Signal_Generate - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;

entity Signal_Generate is
port (

       clk :in  std_logic;
      --Voie de saida c
  
      --Tipo de sinal Type_Wave_Out1 Type_Wave_Out1  P
      
      ---Possibilité de 7 signal 2^3 -1=7 ,  3 bit
       Type_Wave_Out1: in std_logic_vector(2 downto 0):=(others => '0') ;--[sinus=1,square=2]
       Type_Wave_Out2: in std_logic_vector(2 downto 0):=(others => '0');
       ----Gating sont 1->0% , 2->5% , 3->10%,4->15,5->20%,6->50%
       GATING: in std_logic_vector(2 downto 0):=(others => '0');
       ----SORTIE DE 14BIT-----
       OUT1: out std_logic_vector(13 downto 0):=(others => '0') ;
       OUT2: out std_logic_vector(13 downto 0):=(others => '0') 
       );
end Signal_Generate;

architecture Behavioral of Signal_Generate is
signal i : integer range 0 to 2000:=0;
signal U14_SINUS : UNSIGNED(13 downto 0):=(others => '0');

signal U14_SQUARE: UNSIGNED(13 downto 0):=(others => '0'); 
--signal signed1 : UNSIGNED(13 downto 0):=(others => '0');
type memory_type is array (0 to 1999) of integer range 0 to 16384;
--type memory_type is array (0 to 29) of integer range -128 to 127;
--ROM for storing the sine values generated by PYTHON.
--sinus de 2000points ET  FS=125MHz alors 62.5kHz

signal DATA_sinus: memory_type :=(8192,8243,8295,8346,8398,8449,8501,8552,8604,8655,8706,8758,8809,8860,8912,8963,9014,9065,9116,9167,9218,9270
,9321,9371,9422,9473,9524,9575,9625,9676,9727,9777,9828,9878,9928,9979,10029,10079,10129,10179,10229,10279,10328,10378,10427,10477,10526,10576,10625,10674,10723,10772,10821,10869,10918,10966,11015,11063,11111,11159,11207,11255,11302,11350,11397,11445,11492,11539,11586,11633,11679,11726,11772,11818,11864,11910,11956,12002,12047,12092,12138,12183,12227,12272,12317,12361,12405,12449,12493,12537,12580,12624,12667,12710,12753,12795,12838,12880,12922,12964,13006,
13047,13089,13130,13171,13212,13252,13293,13333,13373,13413,13452,13491,13531,13569,13608,13647,13685,13723,13761,13798,13836,13873,13910,13947,13983,14019,14056,14091,14127,14162,14197,14232,14267,14301,14335,14369,14403,14436,14470,14503,14535,14568,14600,14632,14663,14695,14726,14757,14787,14818,14848,14878,14907,14937,14966,14995,15023,15051,15079,15107,15134,15162,15189,15215,15241,15268,15293,15319,15344,15369,15394,15418,15442,15466,15489,15513,15535,15558,15580,15603,15624,15646,15667,15688,15708,15729,15749,15768,15788,15807,15826,15844,15862,15880,15898,15915,15932,15949,15965,15981,15997,16012,16027,16042,16057,16071,16085,16098,16112,16125,16137,16150,16162,16173,16185,16196,16207,16217,16227,16237,16246,16256,16264,16273,16281,16289,16297,16304,16311,16317,16324,16330,16335,16341,16346,16350
,16355,16359,16362,16366,16369,16372,16374,16376,16378,16379,16381,16381,16382,16382,16382,16381,16381,16379,16378,16376,16374,16372,16369,16366,16362,16359,16355,16350,16346,16341,16335,16330,16324,16317,16311,16304,
16297,16289,16281,16273,16264,16256,16246,16237,16227,16217,16207,16196,16185,16173,16162,16150,16137,16125,16112,16098,16085,16071,16057,16042,16027,16012,15997,15981,15965,15949,15932,15915,15898,15880,15862,15844,15826,15807,15788,15768,15749,15729,15708,15688,15667,15646,15624,15603,15580,15558,15535,15513,15489,15466,15442,15418,15394,
15369,15344,15319,15293,15268,15241,15215,15189,15162,15134,15107,15079,15051,15023,14995,14966,14937,14907,14878,14848,14818,14787,14757,14726,14695,14663,14632,14600,14568,14535,14503,14470,14436,14403,14369,14335,14301,14267,14232,14197,14162,14127,14091,14056,14019,13983,13947,13910,13873,13836,13798,13761,13723,13685,13647,13608,13569,13531,13491,13452,13413,13373,13333,13293,13252,13212,13171,13130,13089,13047,13006,
12964,12922,12880,12838,12795,12753,12710,12667,12624,12580,12537,12493,12449,12405,12361,12317,12272,12227,12183,12138,12092,12047,12002,11956,11910,11864,11818,11772,11726,11679,11633,11586,11539,11492,11445,11397,11350,11302,11255,11207,11159,11111,11063,11015,10966,10918,10869,10821,10772,10723,10674,10625,10576,10526,10477,10427,10378,10328,10279,10229,10179,10129,10079,10029,9979,9928,9878,9828,9777,9727,9676,9625,9575,9524,9473,9422,9371,9321,9270,9218,9167,9116,9065,9014,8963,8912,8860,8809,8758,8706,8655,8604,8552,8501,8449,8398,8346,8295,8243,8192,
8141,8089,8038,7986,7935,7883,7832,7780,7729,7678,7626,7575,7524,7472,7421,7370,7319,7268,7217,7166,7114,7063,7013,6962,6911,6860,6809,6759,6708,6657,6607,6556,6506,6456,6405,6355,6305,6255,6205,6155,6105,6056,6006,5957,5907,5858,5808,5759,5710,5661,5612,5563,5515,5466,5418,5369,5321,5273,5225,5177,5129,5082,5034,4987,4939,4892,4845,4798,4751,4705,4658,4612,4566,4520,4474,4428,4382,4337,4292,4246,4201,4157,4112,4067,4023,3979,3935,3891,3847,3804,3760,3717,3674,3631,3589,3546,3504,3462,3420,3378,
3337,3295,3254,3213,3172,3132,3091,3051,3011,2971,2932,2893,2853,2815,2776,2737,2699,2661,2623,2586,2548,2511,2474,2437,2401,2365,2328,2293,2257,2222,2187,2152,2117,2083,2049,2015,1981,1948,1914,1881,1849,1816,1784,1752,1721,1689,1658,1627,1597,1566,1536,1506,1477,1447,1418,1389,1361,1333,1305,1277,1250,1222,1195,1169,1143,1116,1091,1065,1040,1015,990,966,942,918,895,871,849,826,804,781,760,738,717,696,676,655,635,616,596,577,558,540,522,504,486,469,452,435,419,403,
387,372,357,342,327,313,299,286,272,259,247,234,222,211,199,188,177,167,157,147,138,128,120,111,103,95,87,80,73,67,60,54,49,43,38,34,29,25,22,18,15,12,10,8,6,5,3,3,0,0,0,3,3,5,6,8,10,12,15,18,22,25,29,34,38,43,49,54,60,67,73,80,87,95,103,111,120,128,138,147,157,167,177,188,199,211,222,234,247,259,272,286,299,313,327,342,357,372,387,403,419,435,452,469,486,504,522,540,558,577,596,616,635,655,676,696,717,738,760,781,804,826,849,871,895,918,942,966,990,1015,1040,1065,1091,1116,1143,1169,1195,1222,1250,1277,1305,1333,1361,1389,1418,1447,1477,1506,1536,1566,1597,1627,1658,1689,1721,1752,1784,1816,1849,1881,1914,1948,1981,2015,2049,2083,2117,2152,2187,2222,2257,2293,2328,2365,2401,2437,2474,2511,2548,2586,2623,2661,2699,2737,2776,2815,2853,2893,2932,2971,3011,3051,3091,3132,3172,3213,3254,3295,3337,3378,
3420,3462,3504,3546,3589,3631,3674,3717,3760,3804,3847,3891,3935,3979,4023,4067,4112,4157,4201,4246,4292,4337,4382,4428,4474,4520,4566,4612,4658,4705,4751,4798,4845,4892,4939,4987,5034,5082,5129,5177,5225,5273,5321,5369,5418,5466,5515,5563,5612,5661,5710,5759,5808,5858,5907,5957,6006,6056,6105,6155,6205,6255,6305,6355,6405,6456,6506,6556,6607,6657,6708,6759,6809,6860,6911,6962,7013,7063,7114,7166,7217,7268,7319,7370,7421,7472,7524,7575,7626,7678,7729,7780,7832,7883,7935,7986,8038,8089,
8141);


 signal DATA_square0_2000 :memory_type:=(16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
); 
signal DATA_square5_2000 :memory_type:=(16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192
);

signal DATA_square10_2000 :memory_type:=(16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,8192,
8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,8192,
8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192
);

signal DATA_square15_2000 :memory_type:=(
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,
8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,
8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192
);
signal DATA_square20_2000 :memory_type:=(16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192
);
signal DATA_square50_2000 :memory_type:=(
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,8192,
8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,
8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,
8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,
8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,
8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,8192,
8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,
8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,
8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,
8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,
8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192
);
begin

	process(clk)
		begin
			  --to check the rising edge of the clock signal
			if(rising_edge(clk)) then    

				-------------Signal intermediaire -- Passage du DATA en expression de valeur non signe -------------------------------------------
					U14_SINUS <= TO_UNSIGNED(DATA_sinus(i),14);  
					----TRAITEMENT SQUARE CHOIX DE GATING ----
					if(GATING =1)then
					   U14_SQUARE <= TO_UNSIGNED(DATA_square0_2000(i),14);
                    end if ;
                    if(GATING =2)then
					   U14_SQUARE <= TO_UNSIGNED(DATA_square5_2000(i),14);
                    end if ;
                    if(GATING =3)then
					   U14_SQUARE <= TO_UNSIGNED(DATA_square10_2000(i),14);
                    end if ;
                    if(GATING =4)then
					   U14_SQUARE <= TO_UNSIGNED(DATA_square15_2000(i),14);
                    end if ;
                   if(GATING =5)then
					   U14_SQUARE <= TO_UNSIGNED(DATA_square20_2000(i),14);
                    end if ;
                    if(GATING =6)then
					   U14_SQUARE <= TO_UNSIGNED(DATA_square50_2000(i),14);
                    end if ;
                    
					-----------------------Verification et Atribution du type d'onde pour OUT1 ---------------------------------------------------
					if(Type_Wave_Out1 = 1)then
						OUT1<= STD_LOGIC_VECTOR(U14_SINUS); 
					end if;
					if(Type_Wave_Out1 = 2)then
						OUT1<= STD_LOGIC_VECTOR(U14_SQUARE ); 
					end if;

					-----------------------Verification et Atribution du type d'onde pour OUT2 ---------------------------------------------------
					if(Type_Wave_Out2 = 1 )then-- compaison a 1
						OUT2<= STD_LOGIC_VECTOR(U14_SINUS); 
					end if;
					if(Type_Wave_Out2 = 2)then-- compaison a 2
						OUT2<= STD_LOGIC_VECTOR(U14_SQUARE ); 
					end if;


					i <= i+ 1; --INCREMETATION
					if(i = 1999) then
						i <= 0;
					end if;
			end if;
	end process;

end Behavioral;